module imm_gen #(
    REG_WIDTH = 64, INSTRUCTION_WIDTH = 32
) (
    input [INSTRUCTION_WIDTH - 1 : 0] instruction,
    output [REG_WIDTH - 1 : 0] imm 
);
    // finish this module
endmodule